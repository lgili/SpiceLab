* Minimal fallback netlist for PT1000 example
V1 3.3V 0 DC 3.3
R1 3.3V 0 11.3k
.tran 0 1e-3
.end
